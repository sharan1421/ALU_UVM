package alu_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "coverage.sv"
`include "environment.sv"
`include "test.sv"
endpackage
