interface alu_if();
  
  logic [1:0] mode;
  logic [3:0] a;
  logic [3:0] b;
  logic [7:0] y;
  
endinterface:alu_if
